module rvl_ctrl_led_switch_mod # (
  parameter                            RVL_LED_WIDTH       = 8,
  parameter                            RVL_SWITCH_WIDTH    = 8
) (
  input  wire [RVL_LED_WIDTH-1:0]      rvl_leds,
  output wire [RVL_SWITCH_WIDTH-1:0]   rvl_switches
);


endmodule
